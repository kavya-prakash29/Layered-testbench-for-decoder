interface intf();
  
  logic a;
  logic b;
  logic d0;
  logic d1;
  logic d2;
  logic d3;
  
endinterface
